`ifndef _DBB_CHECK_PKG_SVH_
`define _DBB_CHECK_PKG_SVH_
/// UVM DBB CHECK Verification IP Package
   // import uvm_pkg::*;
   // import axi_vip_pkg::*;
   // import axi_vip_dbb_check_pkg::*;
    // DBB transaction
    `include "dbb_check_transaction.sv"            
    // DBB Monitor
    `include "dbb_check_monitor.sv"
    // DBB Scoreboard
    `include "dbb_check_scoreboard.sv"
    // Agents
    `include "dbb_check_agent.sv"

`endif // _DBB_CHECK_PKG_SVH_
